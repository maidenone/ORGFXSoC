`timescale 1 ns/100 ps
// Version: 8.6 8.6.0.34


module eth_pll(POWERDOWN,CLKA,LOCK,GLA);
input POWERDOWN, CLKA;
output  LOCK, GLA;

    wire CLKAP, VCC, GND;
    
    VCC VCC_1_net(.Y(VCC));
    GND GND_1_net(.Y(GND));
    PLL #( .VCOFREQUENCY(125.000) )  Core(.CLKA(CLKAP), .EXTFB(
        GND), .POWERDOWN(POWERDOWN), .GLA(GLA), .LOCK(LOCK), .GLB(
        ), .YB(), .GLC(), .YC(), .OADIV0(GND), .OADIV1(GND), 
        .OADIV2(GND), .OADIV3(GND), .OADIV4(GND), .OAMUX0(GND), 
        .OAMUX1(VCC), .OAMUX2(GND), .DLYGLA0(GND), .DLYGLA1(GND), 
        .DLYGLA2(GND), .DLYGLA3(GND), .DLYGLA4(GND), .OBDIV0(GND), 
        .OBDIV1(GND), .OBDIV2(GND), .OBDIV3(GND), .OBDIV4(GND), 
        .OBMUX0(GND), .OBMUX1(GND), .OBMUX2(GND), .DLYYB0(GND), 
        .DLYYB1(GND), .DLYYB2(GND), .DLYYB3(GND), .DLYYB4(GND), 
        .DLYGLB0(GND), .DLYGLB1(GND), .DLYGLB2(GND), .DLYGLB3(GND)
        , .DLYGLB4(GND), .OCDIV0(GND), .OCDIV1(GND), .OCDIV2(GND), 
        .OCDIV3(GND), .OCDIV4(GND), .OCMUX0(GND), .OCMUX1(GND), 
        .OCMUX2(GND), .DLYYC0(GND), .DLYYC1(GND), .DLYYC2(GND), 
        .DLYYC3(GND), .DLYYC4(GND), .DLYGLC0(GND), .DLYGLC1(GND), 
        .DLYGLC2(GND), .DLYGLC3(GND), .DLYGLC4(GND), .FINDIV0(GND)
        , .FINDIV1(VCC), .FINDIV2(VCC), .FINDIV3(GND), .FINDIV4(
        VCC), .FINDIV5(GND), .FINDIV6(GND), .FBDIV0(GND), .FBDIV1(
        VCC), .FBDIV2(VCC), .FBDIV3(GND), .FBDIV4(VCC), .FBDIV5(
        GND), .FBDIV6(GND), .FBDLY0(GND), .FBDLY1(GND), .FBDLY2(
        GND), .FBDLY3(GND), .FBDLY4(GND), .FBSEL0(VCC), .FBSEL1(
        GND), .XDLYSEL(VCC), .VCOSEL0(GND), .VCOSEL1(GND), 
        .VCOSEL2(VCC));
    PLLINT pllint1(.A(CLKA), .Y(CLKAP));
    
endmodule
